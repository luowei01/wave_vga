// Verilog netlist created by TD v5.0.30786
// Thu Feb 24 19:19:18 2022

`timescale 1ns / 1ps
module wave_ram  // waveram.v(14)
  (
  addra,
  addrb,
  clka,
  clkb,
  dia,
  dib,
  wea,
  web,
  doa,
  dob
  );

  input [9:0] addra;  // waveram.v(37)
  input [9:0] addrb;  // waveram.v(38)
  input clka;  // waveram.v(41)
  input clkb;  // waveram.v(42)
  input [9:0] dia;  // waveram.v(35)
  input [9:0] dib;  // waveram.v(36)
  input wea;  // waveram.v(39)
  input web;  // waveram.v(40)
  output [9:0] doa;  // waveram.v(31)
  output [9:0] dob;  // waveram.v(32)

  parameter ADDR_WIDTH_A = 10;
  parameter ADDR_WIDTH_B = 10;
  parameter DATA_DEPTH_A = 600;
  parameter DATA_DEPTH_B = 600;
  parameter DATA_WIDTH_A = 10;
  parameter DATA_WIDTH_B = 10;
  parameter REGMODE_A = "NOREG";
  parameter REGMODE_B = "NOREG";
  parameter WRITEMODE_A = "NORMAL";
  parameter WRITEMODE_B = "NORMAL";

  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=600;width=9;num_section=1;width_per_section=9;section_size=10;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h00000000000000000000000000000000000000000000000000000000009999B3),
    .INITP_01(256'h70E1E0F81FF000000001FF03E0F0E1C71CE7398CCCE666CCCCD999B333200000),
    .INITP_02(256'h0000000000000000000000000000000000000000003366666CCCE666339CE71C),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h1C1C1C1C1C1C1C1C5C9C4C9C4C8C3C8C3C7C2C7C1C6C1C5C0C5C9C4C9C3C8C2C),
    .INIT_01(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_02(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_03(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_04(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_05(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_06(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_07(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_08(256'h2C7C3C8C3C8C4C9C4C9C5C0C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_09(256'h1C7C2C7C2C8C3C8C4C9C4C0C5C0C6C1C6C2C7C3C8C3C9C4C9C5C0C5C1C6C1C7C),
    .INIT_0A(256'h2C7C1C6C1C5C0C5C0C5C9C4C9C4C9C4C9C4C9C4C9C4C9C5C0C5C0C5C0C6C1C6C),
    .INIT_0B(256'h1C5C8C2C6C9C3C7C0C4C8C2C6C0C4C8C2C6C0C5C9C3C7C2C6C0C5C9C4C8C3C7C),
    .INIT_0C(256'h5C6C8C1C3C5C7C9C2C4C6C9C1C4C6C9C2C5C7C0C3C6C9C2C5C8C1C5C8C1C5C8C),
    .INIT_0D(256'h1C1C1C2C2C2C3C3C4C5C5C6C7C8C9C0C1C2C3C4C5C7C8C9C1C2C4C6C7C9C1C3C),
    .INIT_0E(256'h4C2C1C9C8C7C5C4C3C2C1C0C9C8C7C6C5C5C4C3C3C2C2C2C1C1C1C1C1C1C1C1C),
    .INIT_0F(256'h1C8C5C2C9C6C3C0C7C5C2C9C6C4C1C9C6C4C2C9C7C5C3C0C8C6C4C3C1C9C7C6C),
    .INIT_10(256'h5C0C6C2C7C3C9C4C0C6C2C8C4C0C6C2C8C4C0C7C3C9C6C2C8C5C1C8C5C1C8C5C),
    .INIT_11(256'h0C5C0C4C9C4C9C4C9C4C9C4C9C4C9C4C9C4C0C5C0C5C1C6C1C6C2C7C3C8C4C9C),
    .INIT_12(256'h00000000000000007C2C6C1C6C0C5C0C4C9C4C8C3C8C2C7C2C7C1C6C1C6C0C5C),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_600x10_sub_000000_000 (
    .addra({addra,3'b111}),
    .addrb({addrb,3'b111}),
    .clka(clka),
    .clkb(clkb),
    .dia(dia[8:0]),
    .dib(dib[8:0]),
    .wea(wea),
    .web(web),
    .doa(doa[8:0]),
    .dob(dob[8:0]));
  // address_offset=0;data_offset=9;depth=600;width=1;num_section=1;width_per_section=1;section_size=10;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000010101000000000000000001010101000000010101010000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000010101000000000000000000000000000000000000000000),
    .INIT_09(256'h0000010101010000000001010100000000000000000101010100000001010101),
    .INIT_0A(256'h0000010101010000000000000000000101010100000000010101000000000000),
    .INIT_0B(256'h0101010101010000000000010101010100000000000000000001010101010000),
    .INIT_0C(256'h0101010000000000000000000101010101010100000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000101010101010101),
    .INIT_0E(256'h0101010000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000010101010101010000000000000000000101010101010101),
    .INIT_10(256'h0101000000000000000000010101010100000000000101010101010000000000),
    .INIT_11(256'h0001010100000000010101010000000000000000000101010100000000010101),
    .INIT_12(256'h0000000000000000000000000000010101000000000101010100000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_600x10_sub_000000_009 (
    .addra({addra,3'b111}),
    .addrb({addrb,3'b111}),
    .clka(clka),
    .clkb(clkb),
    .dia({open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,dia[9]}),
    .dib({open_n75,open_n76,open_n77,open_n78,open_n79,open_n80,open_n81,open_n82,dib[9]}),
    .wea(wea),
    .web(web),
    .doa({open_n87,open_n88,open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,doa[9]}),
    .dob({open_n95,open_n96,open_n97,open_n98,open_n99,open_n100,open_n101,open_n102,dob[9]}));

endmodule 

